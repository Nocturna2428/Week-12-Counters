Counter
module counter(btnC,btnU);
  input btnC,btnU;
  output [6:0] data;

